class Packet;
  rand bit [7:0] val;
endclass
