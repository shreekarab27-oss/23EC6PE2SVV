module tb_associative_arrays;

    int mem[int];

endmodule
